package CONSTANTS is
   constant DRCAS : time := 1 ns;
   constant DRCAC : time := 2 ns;
end CONSTANTS;
